`include "./src/sumador/sumador1bPrimitiva.v"

module sumador4b (
    input A, 
    input B, 
    output C,
);
    
endmodule