`include "./src/sumador/sumador1bPrimitiva.v"

module sumador4b (
    input A, 
    input B, 
    output C,
);
    sumador1bPrimitiva s1()
endmodule