`include ""

module alarma_descarga_TB (
);
    reg A;

    initial begin
        
    end
    
endmodule