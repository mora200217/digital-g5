module alarma_descarga (
    ports
);
    
endmodule